module rom_stage_10 (
    input logic         i_clk,
    input logic [8:0]   i_addr,   // [THAY ĐỔI]: 9 bit cho 512 góc
    output logic [31:0] o_data
);

logic [31:0] rom [0:511];

initial begin
    rom[  0] = 32'h00000000; // 0 * -pi/512
    rom[  1] = 32'hfffffe6e; // 1 * -pi/512
    rom[  2] = 32'hfffffcdc; // 2 * -pi/512
    rom[  3] = 32'hfffffb4a; // 3 * -pi/512
    rom[  4] = 32'hfffff9b8; // 4 * -pi/512
    rom[  5] = 32'hfffff825; // 5 * -pi/512
    rom[  6] = 32'hfffff693; // 6 * -pi/512
    rom[  7] = 32'hfffff501; // 7 * -pi/512
    rom[  8] = 32'hfffff36f; // 8 * -pi/512
    rom[  9] = 32'hfffff1dd; // 9 * -pi/512
    rom[ 10] = 32'hfffff04b; // 10 * -pi/512
    rom[ 11] = 32'hffffeeb9; // 11 * -pi/512
    rom[ 12] = 32'hffffed27; // 12 * -pi/512
    rom[ 13] = 32'hffffeb94; // 13 * -pi/512
    rom[ 14] = 32'hffffea02; // 14 * -pi/512
    rom[ 15] = 32'hffffe870; // 15 * -pi/512
    rom[ 16] = 32'hffffe6de; // 16 * -pi/512
    rom[ 17] = 32'hffffe54c; // 17 * -pi/512
    rom[ 18] = 32'hffffe3ba; // 18 * -pi/512
    rom[ 19] = 32'hffffe228; // 19 * -pi/512
    rom[ 20] = 32'hffffe096; // 20 * -pi/512
    rom[ 21] = 32'hffffdf03; // 21 * -pi/512
    rom[ 22] = 32'hffffdd71; // 22 * -pi/512
    rom[ 23] = 32'hffffdbdf; // 23 * -pi/512
    rom[ 24] = 32'hffffda4d; // 24 * -pi/512
    rom[ 25] = 32'hffffd8bb; // 25 * -pi/512
    rom[ 26] = 32'hffffd729; // 26 * -pi/512
    rom[ 27] = 32'hffffd597; // 27 * -pi/512
    rom[ 28] = 32'hffffd405; // 28 * -pi/512
    rom[ 29] = 32'hffffd272; // 29 * -pi/512
    rom[ 30] = 32'hffffd0e0; // 30 * -pi/512
    rom[ 31] = 32'hffffcf4e; // 31 * -pi/512
    rom[ 32] = 32'hffffcdbc; // 32 * -pi/512
    rom[ 33] = 32'hffffcc2a; // 33 * -pi/512
    rom[ 34] = 32'hffffca98; // 34 * -pi/512
    rom[ 35] = 32'hffffc906; // 35 * -pi/512
    rom[ 36] = 32'hffffc774; // 36 * -pi/512
    rom[ 37] = 32'hffffc5e1; // 37 * -pi/512
    rom[ 38] = 32'hffffc44f; // 38 * -pi/512
    rom[ 39] = 32'hffffc2bd; // 39 * -pi/512
    rom[ 40] = 32'hffffc12b; // 40 * -pi/512
    rom[ 41] = 32'hffffbf99; // 41 * -pi/512
    rom[ 42] = 32'hffffbe07; // 42 * -pi/512
    rom[ 43] = 32'hffffbc75; // 43 * -pi/512
    rom[ 44] = 32'hffffbae3; // 44 * -pi/512
    rom[ 45] = 32'hffffb950; // 45 * -pi/512
    rom[ 46] = 32'hffffb7be; // 46 * -pi/512
    rom[ 47] = 32'hffffb62c; // 47 * -pi/512
    rom[ 48] = 32'hffffb49a; // 48 * -pi/512
    rom[ 49] = 32'hffffb308; // 49 * -pi/512
    rom[ 50] = 32'hffffb176; // 50 * -pi/512
    rom[ 51] = 32'hffffafe4; // 51 * -pi/512
    rom[ 52] = 32'hffffae52; // 52 * -pi/512
    rom[ 53] = 32'hffffacbf; // 53 * -pi/512
    rom[ 54] = 32'hffffab2d; // 54 * -pi/512
    rom[ 55] = 32'hffffa99b; // 55 * -pi/512
    rom[ 56] = 32'hffffa809; // 56 * -pi/512
    rom[ 57] = 32'hffffa677; // 57 * -pi/512
    rom[ 58] = 32'hffffa4e5; // 58 * -pi/512
    rom[ 59] = 32'hffffa353; // 59 * -pi/512
    rom[ 60] = 32'hffffa1c1; // 60 * -pi/512
    rom[ 61] = 32'hffffa02e; // 61 * -pi/512
    rom[ 62] = 32'hffff9e9c; // 62 * -pi/512
    rom[ 63] = 32'hffff9d0a; // 63 * -pi/512
    rom[ 64] = 32'hffff9b78; // 64 * -pi/512
    rom[ 65] = 32'hffff99e6; // 65 * -pi/512
    rom[ 66] = 32'hffff9854; // 66 * -pi/512
    rom[ 67] = 32'hffff96c2; // 67 * -pi/512
    rom[ 68] = 32'hffff9530; // 68 * -pi/512
    rom[ 69] = 32'hffff939d; // 69 * -pi/512
    rom[ 70] = 32'hffff920b; // 70 * -pi/512
    rom[ 71] = 32'hffff9079; // 71 * -pi/512
    rom[ 72] = 32'hffff8ee7; // 72 * -pi/512
    rom[ 73] = 32'hffff8d55; // 73 * -pi/512
    rom[ 74] = 32'hffff8bc3; // 74 * -pi/512
    rom[ 75] = 32'hffff8a31; // 75 * -pi/512
    rom[ 76] = 32'hffff889f; // 76 * -pi/512
    rom[ 77] = 32'hffff870c; // 77 * -pi/512
    rom[ 78] = 32'hffff857a; // 78 * -pi/512
    rom[ 79] = 32'hffff83e8; // 79 * -pi/512
    rom[ 80] = 32'hffff8256; // 80 * -pi/512
    rom[ 81] = 32'hffff80c4; // 81 * -pi/512
    rom[ 82] = 32'hffff7f32; // 82 * -pi/512
    rom[ 83] = 32'hffff7da0; // 83 * -pi/512
    rom[ 84] = 32'hffff7c0e; // 84 * -pi/512
    rom[ 85] = 32'hffff7a7b; // 85 * -pi/512
    rom[ 86] = 32'hffff78e9; // 86 * -pi/512
    rom[ 87] = 32'hffff7757; // 87 * -pi/512
    rom[ 88] = 32'hffff75c5; // 88 * -pi/512
    rom[ 89] = 32'hffff7433; // 89 * -pi/512
    rom[ 90] = 32'hffff72a1; // 90 * -pi/512
    rom[ 91] = 32'hffff710f; // 91 * -pi/512
    rom[ 92] = 32'hffff6f7d; // 92 * -pi/512
    rom[ 93] = 32'hffff6dea; // 93 * -pi/512
    rom[ 94] = 32'hffff6c58; // 94 * -pi/512
    rom[ 95] = 32'hffff6ac6; // 95 * -pi/512
    rom[ 96] = 32'hffff6934; // 96 * -pi/512
    rom[ 97] = 32'hffff67a2; // 97 * -pi/512
    rom[ 98] = 32'hffff6610; // 98 * -pi/512
    rom[ 99] = 32'hffff647e; // 99 * -pi/512
    rom[100] = 32'hffff62ec; // 100 * -pi/512
    rom[101] = 32'hffff6159; // 101 * -pi/512
    rom[102] = 32'hffff5fc7; // 102 * -pi/512
    rom[103] = 32'hffff5e35; // 103 * -pi/512
    rom[104] = 32'hffff5ca3; // 104 * -pi/512
    rom[105] = 32'hffff5b11; // 105 * -pi/512
    rom[106] = 32'hffff597f; // 106 * -pi/512
    rom[107] = 32'hffff57ed; // 107 * -pi/512
    rom[108] = 32'hffff565b; // 108 * -pi/512
    rom[109] = 32'hffff54c8; // 109 * -pi/512
    rom[110] = 32'hffff5336; // 110 * -pi/512
    rom[111] = 32'hffff51a4; // 111 * -pi/512
    rom[112] = 32'hffff5012; // 112 * -pi/512
    rom[113] = 32'hffff4e80; // 113 * -pi/512
    rom[114] = 32'hffff4cee; // 114 * -pi/512
    rom[115] = 32'hffff4b5c; // 115 * -pi/512
    rom[116] = 32'hffff49ca; // 116 * -pi/512
    rom[117] = 32'hffff4838; // 117 * -pi/512
    rom[118] = 32'hffff46a5; // 118 * -pi/512
    rom[119] = 32'hffff4513; // 119 * -pi/512
    rom[120] = 32'hffff4381; // 120 * -pi/512
    rom[121] = 32'hffff41ef; // 121 * -pi/512
    rom[122] = 32'hffff405d; // 122 * -pi/512
    rom[123] = 32'hffff3ecb; // 123 * -pi/512
    rom[124] = 32'hffff3d39; // 124 * -pi/512
    rom[125] = 32'hffff3ba7; // 125 * -pi/512
    rom[126] = 32'hffff3a14; // 126 * -pi/512
    rom[127] = 32'hffff3882; // 127 * -pi/512
    rom[128] = 32'hffff36f0; // 128 * -pi/512
    rom[129] = 32'hffff355e; // 129 * -pi/512
    rom[130] = 32'hffff33cc; // 130 * -pi/512
    rom[131] = 32'hffff323a; // 131 * -pi/512
    rom[132] = 32'hffff30a8; // 132 * -pi/512
    rom[133] = 32'hffff2f16; // 133 * -pi/512
    rom[134] = 32'hffff2d83; // 134 * -pi/512
    rom[135] = 32'hffff2bf1; // 135 * -pi/512
    rom[136] = 32'hffff2a5f; // 136 * -pi/512
    rom[137] = 32'hffff28cd; // 137 * -pi/512
    rom[138] = 32'hffff273b; // 138 * -pi/512
    rom[139] = 32'hffff25a9; // 139 * -pi/512
    rom[140] = 32'hffff2417; // 140 * -pi/512
    rom[141] = 32'hffff2285; // 141 * -pi/512
    rom[142] = 32'hffff20f2; // 142 * -pi/512
    rom[143] = 32'hffff1f60; // 143 * -pi/512
    rom[144] = 32'hffff1dce; // 144 * -pi/512
    rom[145] = 32'hffff1c3c; // 145 * -pi/512
    rom[146] = 32'hffff1aaa; // 146 * -pi/512
    rom[147] = 32'hffff1918; // 147 * -pi/512
    rom[148] = 32'hffff1786; // 148 * -pi/512
    rom[149] = 32'hffff15f4; // 149 * -pi/512
    rom[150] = 32'hffff1461; // 150 * -pi/512
    rom[151] = 32'hffff12cf; // 151 * -pi/512
    rom[152] = 32'hffff113d; // 152 * -pi/512
    rom[153] = 32'hffff0fab; // 153 * -pi/512
    rom[154] = 32'hffff0e19; // 154 * -pi/512
    rom[155] = 32'hffff0c87; // 155 * -pi/512
    rom[156] = 32'hffff0af5; // 156 * -pi/512
    rom[157] = 32'hffff0963; // 157 * -pi/512
    rom[158] = 32'hffff07d0; // 158 * -pi/512
    rom[159] = 32'hffff063e; // 159 * -pi/512
    rom[160] = 32'hffff04ac; // 160 * -pi/512
    rom[161] = 32'hffff031a; // 161 * -pi/512
    rom[162] = 32'hffff0188; // 162 * -pi/512
    rom[163] = 32'hfffefff6; // 163 * -pi/512
    rom[164] = 32'hfffefe64; // 164 * -pi/512
    rom[165] = 32'hfffefcd2; // 165 * -pi/512
    rom[166] = 32'hfffefb3f; // 166 * -pi/512
    rom[167] = 32'hfffef9ad; // 167 * -pi/512
    rom[168] = 32'hfffef81b; // 168 * -pi/512
    rom[169] = 32'hfffef689; // 169 * -pi/512
    rom[170] = 32'hfffef4f7; // 170 * -pi/512
    rom[171] = 32'hfffef365; // 171 * -pi/512
    rom[172] = 32'hfffef1d3; // 172 * -pi/512
    rom[173] = 32'hfffef041; // 173 * -pi/512
    rom[174] = 32'hfffeeeae; // 174 * -pi/512
    rom[175] = 32'hfffeed1c; // 175 * -pi/512
    rom[176] = 32'hfffeeb8a; // 176 * -pi/512
    rom[177] = 32'hfffee9f8; // 177 * -pi/512
    rom[178] = 32'hfffee866; // 178 * -pi/512
    rom[179] = 32'hfffee6d4; // 179 * -pi/512
    rom[180] = 32'hfffee542; // 180 * -pi/512
    rom[181] = 32'hfffee3b0; // 181 * -pi/512
    rom[182] = 32'hfffee21d; // 182 * -pi/512
    rom[183] = 32'hfffee08b; // 183 * -pi/512
    rom[184] = 32'hfffedef9; // 184 * -pi/512
    rom[185] = 32'hfffedd67; // 185 * -pi/512
    rom[186] = 32'hfffedbd5; // 186 * -pi/512
    rom[187] = 32'hfffeda43; // 187 * -pi/512
    rom[188] = 32'hfffed8b1; // 188 * -pi/512
    rom[189] = 32'hfffed71f; // 189 * -pi/512
    rom[190] = 32'hfffed58c; // 190 * -pi/512
    rom[191] = 32'hfffed3fa; // 191 * -pi/512
    rom[192] = 32'hfffed268; // 192 * -pi/512
    rom[193] = 32'hfffed0d6; // 193 * -pi/512
    rom[194] = 32'hfffecf44; // 194 * -pi/512
    rom[195] = 32'hfffecdb2; // 195 * -pi/512
    rom[196] = 32'hfffecc20; // 196 * -pi/512
    rom[197] = 32'hfffeca8e; // 197 * -pi/512
    rom[198] = 32'hfffec8fb; // 198 * -pi/512
    rom[199] = 32'hfffec769; // 199 * -pi/512
    rom[200] = 32'hfffec5d7; // 200 * -pi/512
    rom[201] = 32'hfffec445; // 201 * -pi/512
    rom[202] = 32'hfffec2b3; // 202 * -pi/512
    rom[203] = 32'hfffec121; // 203 * -pi/512
    rom[204] = 32'hfffebf8f; // 204 * -pi/512
    rom[205] = 32'hfffebdfd; // 205 * -pi/512
    rom[206] = 32'hfffebc6a; // 206 * -pi/512
    rom[207] = 32'hfffebad8; // 207 * -pi/512
    rom[208] = 32'hfffeb946; // 208 * -pi/512
    rom[209] = 32'hfffeb7b4; // 209 * -pi/512
    rom[210] = 32'hfffeb622; // 210 * -pi/512
    rom[211] = 32'hfffeb490; // 211 * -pi/512
    rom[212] = 32'hfffeb2fe; // 212 * -pi/512
    rom[213] = 32'hfffeb16c; // 213 * -pi/512
    rom[214] = 32'hfffeafd9; // 214 * -pi/512
    rom[215] = 32'hfffeae47; // 215 * -pi/512
    rom[216] = 32'hfffeacb5; // 216 * -pi/512
    rom[217] = 32'hfffeab23; // 217 * -pi/512
    rom[218] = 32'hfffea991; // 218 * -pi/512
    rom[219] = 32'hfffea7ff; // 219 * -pi/512
    rom[220] = 32'hfffea66d; // 220 * -pi/512
    rom[221] = 32'hfffea4db; // 221 * -pi/512
    rom[222] = 32'hfffea349; // 222 * -pi/512
    rom[223] = 32'hfffea1b6; // 223 * -pi/512
    rom[224] = 32'hfffea024; // 224 * -pi/512
    rom[225] = 32'hfffe9e92; // 225 * -pi/512
    rom[226] = 32'hfffe9d00; // 226 * -pi/512
    rom[227] = 32'hfffe9b6e; // 227 * -pi/512
    rom[228] = 32'hfffe99dc; // 228 * -pi/512
    rom[229] = 32'hfffe984a; // 229 * -pi/512
    rom[230] = 32'hfffe96b8; // 230 * -pi/512
    rom[231] = 32'hfffe9525; // 231 * -pi/512
    rom[232] = 32'hfffe9393; // 232 * -pi/512
    rom[233] = 32'hfffe9201; // 233 * -pi/512
    rom[234] = 32'hfffe906f; // 234 * -pi/512
    rom[235] = 32'hfffe8edd; // 235 * -pi/512
    rom[236] = 32'hfffe8d4b; // 236 * -pi/512
    rom[237] = 32'hfffe8bb9; // 237 * -pi/512
    rom[238] = 32'hfffe8a27; // 238 * -pi/512
    rom[239] = 32'hfffe8894; // 239 * -pi/512
    rom[240] = 32'hfffe8702; // 240 * -pi/512
    rom[241] = 32'hfffe8570; // 241 * -pi/512
    rom[242] = 32'hfffe83de; // 242 * -pi/512
    rom[243] = 32'hfffe824c; // 243 * -pi/512
    rom[244] = 32'hfffe80ba; // 244 * -pi/512
    rom[245] = 32'hfffe7f28; // 245 * -pi/512
    rom[246] = 32'hfffe7d96; // 246 * -pi/512
    rom[247] = 32'hfffe7c03; // 247 * -pi/512
    rom[248] = 32'hfffe7a71; // 248 * -pi/512
    rom[249] = 32'hfffe78df; // 249 * -pi/512
    rom[250] = 32'hfffe774d; // 250 * -pi/512
    rom[251] = 32'hfffe75bb; // 251 * -pi/512
    rom[252] = 32'hfffe7429; // 252 * -pi/512
    rom[253] = 32'hfffe7297; // 253 * -pi/512
    rom[254] = 32'hfffe7105; // 254 * -pi/512
    rom[255] = 32'hfffe6f72; // 255 * -pi/512
    rom[256] = 32'hfffe6de0; // 256 * -pi/512
    rom[257] = 32'hfffe6c4e; // 257 * -pi/512
    rom[258] = 32'hfffe6abc; // 258 * -pi/512
    rom[259] = 32'hfffe692a; // 259 * -pi/512
    rom[260] = 32'hfffe6798; // 260 * -pi/512
    rom[261] = 32'hfffe6606; // 261 * -pi/512
    rom[262] = 32'hfffe6474; // 262 * -pi/512
    rom[263] = 32'hfffe62e1; // 263 * -pi/512
    rom[264] = 32'hfffe614f; // 264 * -pi/512
    rom[265] = 32'hfffe5fbd; // 265 * -pi/512
    rom[266] = 32'hfffe5e2b; // 266 * -pi/512
    rom[267] = 32'hfffe5c99; // 267 * -pi/512
    rom[268] = 32'hfffe5b07; // 268 * -pi/512
    rom[269] = 32'hfffe5975; // 269 * -pi/512
    rom[270] = 32'hfffe57e3; // 270 * -pi/512
    rom[271] = 32'hfffe5650; // 271 * -pi/512
    rom[272] = 32'hfffe54be; // 272 * -pi/512
    rom[273] = 32'hfffe532c; // 273 * -pi/512
    rom[274] = 32'hfffe519a; // 274 * -pi/512
    rom[275] = 32'hfffe5008; // 275 * -pi/512
    rom[276] = 32'hfffe4e76; // 276 * -pi/512
    rom[277] = 32'hfffe4ce4; // 277 * -pi/512
    rom[278] = 32'hfffe4b52; // 278 * -pi/512
    rom[279] = 32'hfffe49bf; // 279 * -pi/512
    rom[280] = 32'hfffe482d; // 280 * -pi/512
    rom[281] = 32'hfffe469b; // 281 * -pi/512
    rom[282] = 32'hfffe4509; // 282 * -pi/512
    rom[283] = 32'hfffe4377; // 283 * -pi/512
    rom[284] = 32'hfffe41e5; // 284 * -pi/512
    rom[285] = 32'hfffe4053; // 285 * -pi/512
    rom[286] = 32'hfffe3ec1; // 286 * -pi/512
    rom[287] = 32'hfffe3d2e; // 287 * -pi/512
    rom[288] = 32'hfffe3b9c; // 288 * -pi/512
    rom[289] = 32'hfffe3a0a; // 289 * -pi/512
    rom[290] = 32'hfffe3878; // 290 * -pi/512
    rom[291] = 32'hfffe36e6; // 291 * -pi/512
    rom[292] = 32'hfffe3554; // 292 * -pi/512
    rom[293] = 32'hfffe33c2; // 293 * -pi/512
    rom[294] = 32'hfffe3230; // 294 * -pi/512
    rom[295] = 32'hfffe309d; // 295 * -pi/512
    rom[296] = 32'hfffe2f0b; // 296 * -pi/512
    rom[297] = 32'hfffe2d79; // 297 * -pi/512
    rom[298] = 32'hfffe2be7; // 298 * -pi/512
    rom[299] = 32'hfffe2a55; // 299 * -pi/512
    rom[300] = 32'hfffe28c3; // 300 * -pi/512
    rom[301] = 32'hfffe2731; // 301 * -pi/512
    rom[302] = 32'hfffe259f; // 302 * -pi/512
    rom[303] = 32'hfffe240c; // 303 * -pi/512
    rom[304] = 32'hfffe227a; // 304 * -pi/512
    rom[305] = 32'hfffe20e8; // 305 * -pi/512
    rom[306] = 32'hfffe1f56; // 306 * -pi/512
    rom[307] = 32'hfffe1dc4; // 307 * -pi/512
    rom[308] = 32'hfffe1c32; // 308 * -pi/512
    rom[309] = 32'hfffe1aa0; // 309 * -pi/512
    rom[310] = 32'hfffe190e; // 310 * -pi/512
    rom[311] = 32'hfffe177b; // 311 * -pi/512
    rom[312] = 32'hfffe15e9; // 312 * -pi/512
    rom[313] = 32'hfffe1457; // 313 * -pi/512
    rom[314] = 32'hfffe12c5; // 314 * -pi/512
    rom[315] = 32'hfffe1133; // 315 * -pi/512
    rom[316] = 32'hfffe0fa1; // 316 * -pi/512
    rom[317] = 32'hfffe0e0f; // 317 * -pi/512
    rom[318] = 32'hfffe0c7d; // 318 * -pi/512
    rom[319] = 32'hfffe0aea; // 319 * -pi/512
    rom[320] = 32'hfffe0958; // 320 * -pi/512
    rom[321] = 32'hfffe07c6; // 321 * -pi/512
    rom[322] = 32'hfffe0634; // 322 * -pi/512
    rom[323] = 32'hfffe04a2; // 323 * -pi/512
    rom[324] = 32'hfffe0310; // 324 * -pi/512
    rom[325] = 32'hfffe017e; // 325 * -pi/512
    rom[326] = 32'hfffdffec; // 326 * -pi/512
    rom[327] = 32'hfffdfe59; // 327 * -pi/512
    rom[328] = 32'hfffdfcc7; // 328 * -pi/512
    rom[329] = 32'hfffdfb35; // 329 * -pi/512
    rom[330] = 32'hfffdf9a3; // 330 * -pi/512
    rom[331] = 32'hfffdf811; // 331 * -pi/512
    rom[332] = 32'hfffdf67f; // 332 * -pi/512
    rom[333] = 32'hfffdf4ed; // 333 * -pi/512
    rom[334] = 32'hfffdf35b; // 334 * -pi/512
    rom[335] = 32'hfffdf1c9; // 335 * -pi/512
    rom[336] = 32'hfffdf036; // 336 * -pi/512
    rom[337] = 32'hfffdeea4; // 337 * -pi/512
    rom[338] = 32'hfffded12; // 338 * -pi/512
    rom[339] = 32'hfffdeb80; // 339 * -pi/512
    rom[340] = 32'hfffde9ee; // 340 * -pi/512
    rom[341] = 32'hfffde85c; // 341 * -pi/512
    rom[342] = 32'hfffde6ca; // 342 * -pi/512
    rom[343] = 32'hfffde538; // 343 * -pi/512
    rom[344] = 32'hfffde3a5; // 344 * -pi/512
    rom[345] = 32'hfffde213; // 345 * -pi/512
    rom[346] = 32'hfffde081; // 346 * -pi/512
    rom[347] = 32'hfffddeef; // 347 * -pi/512
    rom[348] = 32'hfffddd5d; // 348 * -pi/512
    rom[349] = 32'hfffddbcb; // 349 * -pi/512
    rom[350] = 32'hfffdda39; // 350 * -pi/512
    rom[351] = 32'hfffdd8a7; // 351 * -pi/512
    rom[352] = 32'hfffdd714; // 352 * -pi/512
    rom[353] = 32'hfffdd582; // 353 * -pi/512
    rom[354] = 32'hfffdd3f0; // 354 * -pi/512
    rom[355] = 32'hfffdd25e; // 355 * -pi/512
    rom[356] = 32'hfffdd0cc; // 356 * -pi/512
    rom[357] = 32'hfffdcf3a; // 357 * -pi/512
    rom[358] = 32'hfffdcda8; // 358 * -pi/512
    rom[359] = 32'hfffdcc16; // 359 * -pi/512
    rom[360] = 32'hfffdca83; // 360 * -pi/512
    rom[361] = 32'hfffdc8f1; // 361 * -pi/512
    rom[362] = 32'hfffdc75f; // 362 * -pi/512
    rom[363] = 32'hfffdc5cd; // 363 * -pi/512
    rom[364] = 32'hfffdc43b; // 364 * -pi/512
    rom[365] = 32'hfffdc2a9; // 365 * -pi/512
    rom[366] = 32'hfffdc117; // 366 * -pi/512
    rom[367] = 32'hfffdbf85; // 367 * -pi/512
    rom[368] = 32'hfffdbdf2; // 368 * -pi/512
    rom[369] = 32'hfffdbc60; // 369 * -pi/512
    rom[370] = 32'hfffdbace; // 370 * -pi/512
    rom[371] = 32'hfffdb93c; // 371 * -pi/512
    rom[372] = 32'hfffdb7aa; // 372 * -pi/512
    rom[373] = 32'hfffdb618; // 373 * -pi/512
    rom[374] = 32'hfffdb486; // 374 * -pi/512
    rom[375] = 32'hfffdb2f4; // 375 * -pi/512
    rom[376] = 32'hfffdb161; // 376 * -pi/512
    rom[377] = 32'hfffdafcf; // 377 * -pi/512
    rom[378] = 32'hfffdae3d; // 378 * -pi/512
    rom[379] = 32'hfffdacab; // 379 * -pi/512
    rom[380] = 32'hfffdab19; // 380 * -pi/512
    rom[381] = 32'hfffda987; // 381 * -pi/512
    rom[382] = 32'hfffda7f5; // 382 * -pi/512
    rom[383] = 32'hfffda663; // 383 * -pi/512
    rom[384] = 32'hfffda4d0; // 384 * -pi/512
    rom[385] = 32'hfffda33e; // 385 * -pi/512
    rom[386] = 32'hfffda1ac; // 386 * -pi/512
    rom[387] = 32'hfffda01a; // 387 * -pi/512
    rom[388] = 32'hfffd9e88; // 388 * -pi/512
    rom[389] = 32'hfffd9cf6; // 389 * -pi/512
    rom[390] = 32'hfffd9b64; // 390 * -pi/512
    rom[391] = 32'hfffd99d2; // 391 * -pi/512
    rom[392] = 32'hfffd983f; // 392 * -pi/512
    rom[393] = 32'hfffd96ad; // 393 * -pi/512
    rom[394] = 32'hfffd951b; // 394 * -pi/512
    rom[395] = 32'hfffd9389; // 395 * -pi/512
    rom[396] = 32'hfffd91f7; // 396 * -pi/512
    rom[397] = 32'hfffd9065; // 397 * -pi/512
    rom[398] = 32'hfffd8ed3; // 398 * -pi/512
    rom[399] = 32'hfffd8d41; // 399 * -pi/512
    rom[400] = 32'hfffd8bae; // 400 * -pi/512
    rom[401] = 32'hfffd8a1c; // 401 * -pi/512
    rom[402] = 32'hfffd888a; // 402 * -pi/512
    rom[403] = 32'hfffd86f8; // 403 * -pi/512
    rom[404] = 32'hfffd8566; // 404 * -pi/512
    rom[405] = 32'hfffd83d4; // 405 * -pi/512
    rom[406] = 32'hfffd8242; // 406 * -pi/512
    rom[407] = 32'hfffd80b0; // 407 * -pi/512
    rom[408] = 32'hfffd7f1d; // 408 * -pi/512
    rom[409] = 32'hfffd7d8b; // 409 * -pi/512
    rom[410] = 32'hfffd7bf9; // 410 * -pi/512
    rom[411] = 32'hfffd7a67; // 411 * -pi/512
    rom[412] = 32'hfffd78d5; // 412 * -pi/512
    rom[413] = 32'hfffd7743; // 413 * -pi/512
    rom[414] = 32'hfffd75b1; // 414 * -pi/512
    rom[415] = 32'hfffd741f; // 415 * -pi/512
    rom[416] = 32'hfffd728c; // 416 * -pi/512
    rom[417] = 32'hfffd70fa; // 417 * -pi/512
    rom[418] = 32'hfffd6f68; // 418 * -pi/512
    rom[419] = 32'hfffd6dd6; // 419 * -pi/512
    rom[420] = 32'hfffd6c44; // 420 * -pi/512
    rom[421] = 32'hfffd6ab2; // 421 * -pi/512
    rom[422] = 32'hfffd6920; // 422 * -pi/512
    rom[423] = 32'hfffd678e; // 423 * -pi/512
    rom[424] = 32'hfffd65fb; // 424 * -pi/512
    rom[425] = 32'hfffd6469; // 425 * -pi/512
    rom[426] = 32'hfffd62d7; // 426 * -pi/512
    rom[427] = 32'hfffd6145; // 427 * -pi/512
    rom[428] = 32'hfffd5fb3; // 428 * -pi/512
    rom[429] = 32'hfffd5e21; // 429 * -pi/512
    rom[430] = 32'hfffd5c8f; // 430 * -pi/512
    rom[431] = 32'hfffd5afd; // 431 * -pi/512
    rom[432] = 32'hfffd596a; // 432 * -pi/512
    rom[433] = 32'hfffd57d8; // 433 * -pi/512
    rom[434] = 32'hfffd5646; // 434 * -pi/512
    rom[435] = 32'hfffd54b4; // 435 * -pi/512
    rom[436] = 32'hfffd5322; // 436 * -pi/512
    rom[437] = 32'hfffd5190; // 437 * -pi/512
    rom[438] = 32'hfffd4ffe; // 438 * -pi/512
    rom[439] = 32'hfffd4e6c; // 439 * -pi/512
    rom[440] = 32'hfffd4cda; // 440 * -pi/512
    rom[441] = 32'hfffd4b47; // 441 * -pi/512
    rom[442] = 32'hfffd49b5; // 442 * -pi/512
    rom[443] = 32'hfffd4823; // 443 * -pi/512
    rom[444] = 32'hfffd4691; // 444 * -pi/512
    rom[445] = 32'hfffd44ff; // 445 * -pi/512
    rom[446] = 32'hfffd436d; // 446 * -pi/512
    rom[447] = 32'hfffd41db; // 447 * -pi/512
    rom[448] = 32'hfffd4049; // 448 * -pi/512
    rom[449] = 32'hfffd3eb6; // 449 * -pi/512
    rom[450] = 32'hfffd3d24; // 450 * -pi/512
    rom[451] = 32'hfffd3b92; // 451 * -pi/512
    rom[452] = 32'hfffd3a00; // 452 * -pi/512
    rom[453] = 32'hfffd386e; // 453 * -pi/512
    rom[454] = 32'hfffd36dc; // 454 * -pi/512
    rom[455] = 32'hfffd354a; // 455 * -pi/512
    rom[456] = 32'hfffd33b8; // 456 * -pi/512
    rom[457] = 32'hfffd3225; // 457 * -pi/512
    rom[458] = 32'hfffd3093; // 458 * -pi/512
    rom[459] = 32'hfffd2f01; // 459 * -pi/512
    rom[460] = 32'hfffd2d6f; // 460 * -pi/512
    rom[461] = 32'hfffd2bdd; // 461 * -pi/512
    rom[462] = 32'hfffd2a4b; // 462 * -pi/512
    rom[463] = 32'hfffd28b9; // 463 * -pi/512
    rom[464] = 32'hfffd2727; // 464 * -pi/512
    rom[465] = 32'hfffd2594; // 465 * -pi/512
    rom[466] = 32'hfffd2402; // 466 * -pi/512
    rom[467] = 32'hfffd2270; // 467 * -pi/512
    rom[468] = 32'hfffd20de; // 468 * -pi/512
    rom[469] = 32'hfffd1f4c; // 469 * -pi/512
    rom[470] = 32'hfffd1dba; // 470 * -pi/512
    rom[471] = 32'hfffd1c28; // 471 * -pi/512
    rom[472] = 32'hfffd1a96; // 472 * -pi/512
    rom[473] = 32'hfffd1903; // 473 * -pi/512
    rom[474] = 32'hfffd1771; // 474 * -pi/512
    rom[475] = 32'hfffd15df; // 475 * -pi/512
    rom[476] = 32'hfffd144d; // 476 * -pi/512
    rom[477] = 32'hfffd12bb; // 477 * -pi/512
    rom[478] = 32'hfffd1129; // 478 * -pi/512
    rom[479] = 32'hfffd0f97; // 479 * -pi/512
    rom[480] = 32'hfffd0e05; // 480 * -pi/512
    rom[481] = 32'hfffd0c72; // 481 * -pi/512
    rom[482] = 32'hfffd0ae0; // 482 * -pi/512
    rom[483] = 32'hfffd094e; // 483 * -pi/512
    rom[484] = 32'hfffd07bc; // 484 * -pi/512
    rom[485] = 32'hfffd062a; // 485 * -pi/512
    rom[486] = 32'hfffd0498; // 486 * -pi/512
    rom[487] = 32'hfffd0306; // 487 * -pi/512
    rom[488] = 32'hfffd0174; // 488 * -pi/512
    rom[489] = 32'hfffcffe1; // 489 * -pi/512
    rom[490] = 32'hfffcfe4f; // 490 * -pi/512
    rom[491] = 32'hfffcfcbd; // 491 * -pi/512
    rom[492] = 32'hfffcfb2b; // 492 * -pi/512
    rom[493] = 32'hfffcf999; // 493 * -pi/512
    rom[494] = 32'hfffcf807; // 494 * -pi/512
    rom[495] = 32'hfffcf675; // 495 * -pi/512
    rom[496] = 32'hfffcf4e3; // 496 * -pi/512
    rom[497] = 32'hfffcf350; // 497 * -pi/512
    rom[498] = 32'hfffcf1be; // 498 * -pi/512
    rom[499] = 32'hfffcf02c; // 499 * -pi/512
    rom[500] = 32'hfffcee9a; // 500 * -pi/512
    rom[501] = 32'hfffced08; // 501 * -pi/512
    rom[502] = 32'hfffceb76; // 502 * -pi/512
    rom[503] = 32'hfffce9e4; // 503 * -pi/512
    rom[504] = 32'hfffce852; // 504 * -pi/512
    rom[505] = 32'hfffce6bf; // 505 * -pi/512
    rom[506] = 32'hfffce52d; // 506 * -pi/512
    rom[507] = 32'hfffce39b; // 507 * -pi/512
    rom[508] = 32'hfffce209; // 508 * -pi/512
    rom[509] = 32'hfffce077; // 509 * -pi/512
    rom[510] = 32'hfffcdee5; // 510 * -pi/512
    rom[511] = 32'hfffcdd53; // 511 * -pi/512
end

always @(posedge i_clk) begin
    o_data <= rom[i_addr];
end

endmodule
