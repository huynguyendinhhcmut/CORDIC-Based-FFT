module stage_1 (	
	input logic i_clk, i_reset
);

endmodule